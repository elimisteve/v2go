module main

println('Hello, World!')
